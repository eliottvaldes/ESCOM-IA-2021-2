library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity adder4b is
PORT(
A,B:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
S:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
CI:IN STD_LOGIC;
C0:OUT STD_LOGIC);
end adder4b;
architecture Behavioral of adder4b is
SIGNAL SC:STD_LOGIC_VECTOR(3 DOWNTO 0);
COMPONENT FullADDER
PORT(
CI,A,B:IN STD_LOGIC;
S,C0:OUT STD_LOGIC);
END COMPONENT;
begin
U0:FullADDER
PORT MAP(CI,A(0),B(0),S(0),SC(0));
U1_U3:
FOR I IN 1 TO 2 GENERATE
U:FullADDER PORT MAP(SC(I-1),A(I),B(I),S(I),SC(I));
END GENERATE;
U4:FullADDER PORT MAP(SC(2),A(3),B(3),S(3),C0);
end Behavioral;
